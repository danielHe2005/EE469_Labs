// Test bench for Register file
`timescale 1ns/10ps

module regstim(); 		

	parameter ClockDelay = 5000;

	logic	[4:0] 	ReadRegister1, ReadRegister2, WriteRegister;
	logic [63:0]	WriteData;
	logic 			RegWrite, clk;
	logic [63:0]	ReadData1, ReadData2;

	integer i;

	// Your register file MUST be named "regfile".
	// Also you must make sure that the port declarations
	// match up with the module instance in this stimulus file.
	regfile dut (.ReadData1, .ReadData2, .WriteData, 
					 .ReadRegister1, .ReadRegister2, .WriteRegister,
					 .RegWrite, .clk);

	// Force %t's to print in a nice format.
	initial $timeformat(-9, 2, " ns", 10);

	initial begin // Set up the clock
		clk <= 0;
		forever #(ClockDelay/2) clk <= ~clk;
	end

	initial begin
		// Try to write the value 0xA0 into register 31.
		// Register 31 should always be at the value of 0.
		RegWrite <= 5'd0;
		ReadRegister1 <= 5'd31;
		ReadRegister2 <= 5'd0;
		WriteRegister <= 5'd31;
		WriteData <= 64'h00000000000000A0;
		@(posedge clk);
		
		$display("%t Attempting overwrite of register 31, which should always be 0", $time);
		RegWrite <= 1;
		@(posedge clk);
		$display("WriteData=%0d, out=%0d (expected %0d)", WriteData, ReadData1, 64'd0); // creates a display to show the intended and actual results of attempting to overwrite Register 31
      assert (ReadData1 == 64'd0) else $error("Register 31 was overwritten to %0d, test failed", ReadData1);

		// Write a value into each  register.
		$display("%t Writing pattern to all registers.", $time);
		for (i=0; i<31; i=i+1) begin
			RegWrite <= 0;
			ReadRegister1 <= i-1;
			ReadRegister2 <= i;
			WriteRegister <= i;
			WriteData <= i*64'h0000010204080001;
			@(posedge clk);
			$display("WriteData=%0d, out=%0d", WriteData, ReadData2); // creates a display to show that the write value hasn't been written into the designated write register yet
			assert ($isunknown(ReadData2)) else $error("Register %0d has been overwritten to %0d even though RegWrite was false, test failed", i, ReadData2);
			RegWrite <= 1;
			@(posedge clk);
			@(posedge clk);
			$display("WriteData=%0d, out=%0d (expected %0d)", WriteData, ReadData2, WriteData); // creates a display to show that the write value is now written to the designated write register
			assert (ReadData2 == WriteData) else $error("Register %0d was not written to %0d, test failed", i, WriteData);
		end

		// Go back and verify that the registers
		// retained the data.
		$display("%t Checking pattern.", $time);
		for (i=0; i<32; i=i+1) begin
			RegWrite <= 0;
			ReadRegister1 <= i-1;
			ReadRegister2 <= i;
			WriteRegister <= i;
			WriteData <= i*64'h0000000000000100+i;
			@(posedge clk);
		end
		$stop;
	end
endmodule